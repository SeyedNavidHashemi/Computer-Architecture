`timescale 1ns/1ns

module divider(AIN , BIN , START , SCLR , CLK , QOUT , DVZ , OVF , BUSY , VALID);
    input [9:0] AIN , BIN;
    input START , SCLR , CLK;
    output [9:0] QOUT;
    output DVZ , OVF , BUSY , VALID;
    wire DEC_CNT, LD_CNT, SEL_CNT, LD_A, LD_B, LD_ACC, SH_ACC, LD_Q, SH_Q, SET_F, RESET_F, SEL_X, AGTB_CNT , ALL_ZERO, AGTB, B_IS_ZERO, COUT, SET_NEW, RESET_NEW, FINISHORNOT;
    
    datapath dp(AIN, BIN, DEC_CNT, LD_CNT, SEL_CNT, CLK, SCLR, LD_A, LD_B, LD_ACC, SH_ACC, LD_Q, SH_Q, SET_F, RESET_F, SEL_X, QOUT, ALL_ZERO, AGTB, B_IS_ZERO, COUT, SET_NEW, RESET_NEW, FINISHORNOT);

    controller cu(START, CLK, SCLR, AGTB, ALL_ZERO, B_IS_ZERO, COUT, LD_A, LD_B, LD_ACC, SH_ACC, LD_Q, SH_Q, SEL_X, SET_F, RESET_F, SET_NEW, RESET_NEW, FINISHORNOT, OVF, VALID, BUSY, DVZ, DEC_CNT, LD_CNT, SEL_CNT);
endmodule